netcdf s3__sy_2_syrtax {
dimensions:
	AMIN = 40 ;
	ADA = 31 ;
	SZA = 20 ;
	OLC_VZA = 18 ;
	SLN_VZA = 18 ;
	SLO_VZA = 1 ;
	air_pressure = 4 ;
	water_vapour = 3 ;
	T550 = 11 ;
	OLC_channel = 18 ;
	SLN_channel = 6 ;
	SLO_channel = 6 ;
	SYN_channel = 30 ;
	SLS_band = 6 ;
variables:
	float ADA(ADA) ;
		ADA:long_name = "Azimuth difference angle" ;
		ADA:units = "degrees" ;
		ADA:valid_min = 0.f ;
		ADA:valid_max = 180.f ;
	float SZA(SZA) ;
		SZA:long_name = "Solar zenith angle" ;
		SZA:units = "degrees" ;
		SZA:valid_min = 0.f ;
		SZA:valid_max = 70.f ;
		SZA:standard_name = "solar_zenith_angle" ;
	float OLC_VZA(OLC_VZA) ;
		OLC_VZA:long_name = "OLCI view zenith angle" ;
		OLC_VZA:valid_min = 0.f ;
		OLC_VZA:valid_max = 55.f ;
	float SLN_VZA(SLN_VZA) ;
		SLN_VZA:long_name = "SLSTR nadir view zenith angle" ;
		SLN_VZA:units = "degrees" ;
		SLN_VZA:valid_min = 6.f ;
		SLN_VZA:valid_max = 58.f ;
	float SLO_VZA(SLO_VZA) ;
		SLO_VZA:long_name = "SLSTR oblique view zenith angle" ;
		SLO_VZA:units = "degrees" ;
		SLO_VZA:valid_min = 55.f ;
		SLO_VZA:valid_max = 55.f ;
	float air_pressure(air_pressure) ;
		air_pressure:long_name = "Surface pressure" ;
		air_pressure:units = "hPa" ;
		air_pressure:valid_min = 800.f ;
		air_pressure:valid_max = 1030.f ;
		air_pressure:standard_name = "air_pressure_at_sea_level" ;
	float water_vapour(water_vapour) ;
		water_vapour:long_name = "Total column water vapour" ;
		water_vapour:units = "g cm-2" ;
		water_vapour:valid_min = 0.f ;
		water_vapour:valid_max = 5.f ;
	short AMIN(AMIN) ;
		AMIN:long_name = "Aerosol model index number" ;
		AMIN:valid_min = 1 ;
		AMIN:valid_max = 40 ;
	float T550(T550) ;
		T550:long_name = "Aerosol optical thickness" ;
		T550:valid_min = 0.f ;
		T550:valid_max = 4.f ;
		T550:standard_name = "atmosphere_optical_thickness_due_to_aerosol" ;
	short OLC_channel(OLC_channel) ;
		OLC_channel:long_name = "SYN channel index number" ;
		OLC_channel:valid_min = 1 ;
		OLC_channel:valid_max = 18 ;
	short SLN_channel(SLN_channel) ;
		SLN_channel:long_name = "SYN channel index number" ;
		SLN_channel:valid_min = 19 ;
		SLN_channel:valid_max = 24 ;
	short SLO_channel(SLO_channel) ;
		SLO_channel:long_name = "SYN channel index number" ;
		SLO_channel:valid_min = 25 ;
		SLO_channel:valid_max = 30 ;
	short SYN_channel(SYN_channel) ;
		SYN_channel:long_name = "SYN channel index number" ;
		SYN_channel:valid_min = 1 ;
		SYN_channel:valid_max = 30 ;
	short SLS_band(SLS_band) ;
		SLS_band:valid_min = 1 ;
		SLS_band:valid_max = 6 ;
	ubyte OLC_R_atm(ADA, SZA, OLC_VZA, air_pressure, water_vapour, T550, AMIN, OLC_channel) ;
		OLC_R_atm:long_name = "Atmospheric scattering term" ;
		OLC_R_atm:scale_factor = 0.004;
		OLC_R_atm:valid_min = 0u ;
		OLC_R_atm:valid_max = 250u ;
	ubyte SLN_R_atm(ADA, SZA, SLN_VZA, air_pressure, water_vapour, T550, AMIN, SLN_channel) ;
		SLN_R_atm:long_name = "Atmospheric scattering term" ;
		SLN_R_atm:scale_factor = 0.004;
		SLN_R_atm:valid_min = 0 ;
		SLN_R_atm:valid_max = 250 ;
	ubyte SLO_R_atm(ADA, SZA, SLO_VZA, air_pressure, water_vapour, T550, AMIN, SLO_channel) ;
		SLO_R_atm:long_name = "Atmospheric scattering term" ;
		SLO_R_atm:scale_factor = 0.004;
		SLO_R_atm:valid_min = 0 ;
		SLO_R_atm:valid_max = 250 ;
	float t(SZA, air_pressure, water_vapour, T550, AMIN, SYN_channel) ;
		t:long_name = "Atmospheric transmission" ;
		t:valid_min = 0.0 ;
		t:valid_max = 1.0 ;
	float rho_atm(air_pressure, water_vapour, T550, AMIN, SYN_channel) ;
		rho_atm:long_name = "Atmospheric bihemispherical Albedo" ;
		rho_atm:valid_min = 0.0 ;
		rho_atm:valid_max = 1.0 ;
	float D(SZA, air_pressure, T550, AMIN, SLS_band) ;
		D:long_name = "Fraction of diffuse irradiance" ;
		D:valid_min = 0.0 ;
		D:valid_max = 1.0 ;
	float C_O3(SYN_channel) ;
		C_O3:long_name = "Ozone correction factor" ;
		C_O3:valid_min = 0.0 ;
		C_O3:valid_max = 1.0 ;
	float A550(AMIN) ;
		A550:standard_name = "aerosol_angstrom_exponent" ;
		A550:valid_min = -0.5 ;
		A550:valid_max = 2.5 ;
	float delta_rt ;
		delta_rt:valid_min = 0.0 ;
		delta_rt:valid_max = 1.0 ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "SYN L2 radiative transfer simulation dataset" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-L2-SD-08-S-BC-IODD" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "S3__SY_2_SYRTAX_20110701T000000_20120701T000000_20112007T120000__BC__D_NT_AUX_01.nc" ;
		:creation_time = "20110720T120000Z" ;
		:validity_start = "20110701T000000Z" ;
		:validity_stop = "20120701T000000Z" ;
data:

 ADA = 0.f, 6.f, 12.f, 18.f, 24.f, 30.f, 36.f, 42.f, 48.f, 54.f, 60.f, 66.f, 72.f, 78.f, 84.f, 90.f, 96.f, 102.f,
    108.f, 114.f, 120.f, 126.f, 132.f, 138.f, 144.f, 150.f, 156.f, 162.f, 168.f, 174.f, 180.f ;

 SZA = 0.f, 3.5f, 7.f, 11.5f, 14.f, 17.5f, 21.f, 24.5f, 28.f, 31.5f, 34.f, 37.5f, 41.f, 44.5f, 48.f, 51.5f, 54.f,
    57.5f, 61.f, 70.f ;

 OLC_VZA = 0.0f, 3.0f, 6.0f, 9.0f, 12.0f, 15.0f, 18.0f, 21.0f, 24.0f, 27.0f, 30.0f, 33.0f, 36.0f, 39.0f, 42.0f, 45.0f, 50.0f, 55.0f ;

 SLN_VZA = 6.0f, 9.0f, 12.0f, 15.0f, 18.0f, 21.0f, 24.0f, 27.0f, 30.0f, 33.0f, 36.0f, 39.0f, 42.0f, 45.0f, 48.0f, 51.0f, 54.0f, 58.0f ;

 SLO_VZA = 55.0f ;

 air_pressure = 800.f, 900.f, 1000.f, 1030.f ;

 water_vapour = 0.f, 2.f, 5.f ;

 AMIN = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23,
    24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

 T550 = 0.f, 0.05f, 0.1f, 0.2f, 0.4f, 0.6f, 1.f, 1.5f, 2.f, 3.f, 4.f ;

 OLC_channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18 ;

 SLN_channel = 19, 20, 21, 22, 23, 24 ;

 SLO_channel = 25, 26, 27, 28, 29, 30 ;

 SYN_channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30 ;

 SLS_band = 1, 2, 3, 4, 5, 6 ;

 OLC_R_atm = ${OLC_R_ATM} ;

 SLN_R_atm = ${SLN_R_ATM} ;

 SLO_R_atm = ${SLO_R_ATM} ;

 t  = ${T} ;

 rho_atm  = ${RHO_ATM} ;

 D =  ${D} ;

 C_O3 =  0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f, 0.f,
    0.f, 0.f, 0.f, 0.f, 0.f 0.f,
    0.f, 0.f, 0.f, 0.f, 0.f 0.f ;

 delta_rt = 0.005f;
}
