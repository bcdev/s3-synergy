netcdf s3__sy_2_syrtax {
dimensions:
	AMIN = 40 ;
	ADA = 31 ;
	SZA = 20 ;
	OLC_VZA = 18 ;
	SLN_VZA = 18 ;
	SLO_VZA = 1 ;
	air_pressure = 4 ;
	water_vapour = 3 ;
	T550 = 11 ;
	OLC_channel = 18 ;
	SLN_channel = 6 ;
	SLO_channel = 6 ;
	SYN_channel = 30 ;
	SLS_band = 6 ;
variables:
	float ADA(ADA) ;
		ADA:long_name = "Azimuth difference angle" ;
		ADA:units = "degrees" ;
		ADA:valid_min = 0.f ;
		ADA:valid_max = 180.f ;
	float SZA(SZA) ;
		SZA:long_name = "Solar zenith angle" ;
		SZA:units = "degrees" ;
		SZA:valid_min = 0.f ;
		SZA:valid_max = 70.f ;
		SZA:standard_name = "solar_zenith_angle" ;
	float OLC_VZA(OLC_VZA) ;
		OLC_VZA:long_name = "OLCI view zenith angle" ;
		OLC_VZA:valid_min = 0.f ;
		OLC_VZA:valid_max = 55.f ;
	float SLN_VZA(SLN_VZA) ;
		SLN_VZA:long_name = "SLSTR nadir view zenith angle" ;
		SLN_VZA:units = "degrees" ;
		SLN_VZA:valid_min = 6.f ;
		SLN_VZA:valid_max = 58.f ;
	float SLO_VZA(SLO_VZA) ;
		SLO_VZA:long_name = "SLSTR oblique view zenith angle" ;
		SLO_VZA:units = "degrees" ;
		SLO_VZA:valid_min = 55.f ;
		SLO_VZA:valid_max = 55.f ;
	float air_pressure(air_pressure) ;
		air_pressure:long_name = "Surface pressure" ;
		air_pressure:units = "hPa" ;
		air_pressure:valid_min = 800.f ;
		air_pressure:valid_max = 1030.f ;
		air_pressure:standard_name = "air_pressure_at_sea_level" ;
	float water_vapour(water_vapour) ;
		water_vapour:long_name = "Total column water vapour" ;
		water_vapour:units = "g cm-2" ;
		water_vapour:valid_min = 0.f ;
		water_vapour:valid_max = 5.f ;
	short AMIN(AMIN) ;
		AMIN:long_name = "Aerosol model index number" ;
		AMIN:valid_min = 1 ;
		AMIN:valid_max = 40 ;
	float T550(T550) ;
		T550:long_name = "Aerosol optical thickness" ;
		T550:valid_min = 0.f ;
		T550:valid_max = 4.f ;
		T550:standard_name = "atmosphere_optical_thickness_due_to_aerosol" ;
	short OLC_channel(OLC_channel) ;
		OLC_channel:long_name = "SYN channel index number" ;
		OLC_channel:valid_min = 1.f ;
		OLC_channel:valid_max = 18.f ;
	short SLN_channel(SLN_channel) ;
		SLN_channel:long_name = "SYN channel index number" ;
		SLN_channel:valid_min = 19.f ;
		SLN_channel:valid_max = 24.f ;
	short SLO_channel(SLO_channel) ;
		SLO_channel:long_name = "SYN channel index number" ;
		SLO_channel:valid_min = 25.f ;
		SLO_channel:valid_max = 30.f ;
	short SYN_channel(SYN_channel) ;
		SYN_channel:long_name = "SYN channel index number" ;
		SYN_channel:valid_min = 1.f ;
		SYN_channel:valid_max = 30.f ;
	short SLS_band(SLS_band) ;
		SLS_band:valid_min = 1 ;
		SLS_band:valid_max = 6 ;
	ubyte OLC_R_atm(ADA, SZA, OLC_VZA, air_pressure, water_vapour, T550, AMIN, OLC_channel) ;
		OLC_R_atm:long_name = "Atmospheric scattering term" ;
		OLC_R_atm:scale_factor = 0.004;
		OLC_R_atm:valid_min = 0 ;
		OLC_R_atm:valid_max = 250 ;
	ubyte SLN_R_atm(ADA, SZA, SLN_VZA, air_pressure, water_vapour, T550, AMIN, SLN_channel) ;
		SLN_R_atm:long_name = "Atmospheric scattering term" ;
		SLN_R_atm:scale_factor = 0.004;
		SLN_R_atm:valid_min = 0 ;
		SLN_R_atm:valid_max = 250 ;
	ubyte SLO_R_atm(ADA, SZA, SLO_VZA, air_pressure, water_vapour, T550, AMIN, SLO_channel) ;
		SLO_R_atm:long_name = "Atmospheric scattering term" ;
		SLO_R_atm:scale_factor = 0.004;
		SLO_R_atm:valid_min = 0 ;
		SLO_R_atm:valid_max = 250 ;
	float t(SZA, air_pressure, water_vapour, T550, AMIN, SYN_channel) ;
		t:long_name = "Atmospheric transmission" ;
		t:valid_min = 0.0 ;
		t:valid_max = 1.0 ;
	float rho_atm(air_pressure, water_vapour, T550, AMIN, SYN_channel) ;
		rho_atm:long_name = "Atmospheric bihemispherical Albedo" ;
		rho_atm:valid_min = 0.0 ;
		rho_atm:valid_max = 1.0 ;
	float D(SZA, air_pressure, T550, AMIN, SLS_band) ;
		D:long_name = "Fraction of diffuse irradiance" ;
		D:valid_min = 0.0 ;
		D:valid_max = 1.0 ;
	float C_O3(SYN_channel) ;
		C_O3:long_name = "Ozone correction factor" ;
		C_O3:valid_min = 0.0 ;
		C_O3:valid_max = 1.0 ;
	float A550(AMIN) ;
		A550:standard_name = "aerosol_angstrom_exponent" ;
		A550:valid_min = -0.5 ;
		A550:valid_max = 2.5 ;
	float delta_rt ;
		delta_rt:valid_min = 0.0 ;
		delta_rt:valid_max = 1.0 ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "SYN L2 radiative transfer simulation dataset" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-L2-SD-08-S-BC-IODD" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "S3__SY_2_SYRTAX_20101201T000000_20110301T000000_20101207T120000__BC__D_NT_AUX_01.nc" ;
		:creation_time = "20101207T120000Z" ;
		:validity_start = "20101201T000000Z" ;
		:validity_stop = "20110301T000000Z" ;
data:

 ADA = 0, 6, 12, 18, 24, 30, 36, 42, 48, 54, 60, 66, 72, 78, 84, 90, 96, 102, 
    108, 114, 120, 126, 132, 138, 144, 150, 156, 162, 168, 174, 180 ;

 SZA = -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, -1, 
    -1, -1, -1 ;

 OLC_VZA = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SLN_VZA = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 SLO_VZA = _ ;

 air_pressure = 800, 900, 1000, 1030 ;

 water_vapour = 0, 2, 5 ;

 AMIN = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _ ;

 T550 = 0, 0.05, 0.1, 0.2, 0.4, 0.6, 1, 1.5, 2, 3, 4 ;

 OLC_channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18 ;

 SLN_channel = 19, 20, 21, 22, 23, 24 ;

 SLO_channel = 25, 26, 27, 28, 29, 30 ;

 SYN_channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30 ;

 delta_rt = 0.005;
}