netcdf s3__sy_2_vsrtax {
dimensions:
	AMIN = 40 ;
	ADA = 31 ;
	SZA = 20 ;
	VZA = 18 ;
	air_pressure = 4 ;
	water_vapour = 3 ;
	T550 = 11 ;
	channel = 4;
variables:
	float ADA(ADA) ;
		ADA:long_name = "Azimuth difference angle" ;
		ADA:units = "degrees" ;
		ADA:valid_min = 0.f ;
		ADA:valid_max = 180.f ;
	float SZA(SZA) ;
		SZA:long_name = "Solar zenith angle" ;
		SZA:units = "degrees" ;
		SZA:valid_min = 0.f ;
		SZA:valid_max = 70.f ;
		SZA:standard_name = "solar_zenith_angle" ;
	float VZA(VZA) ;
		VZA:long_name = "View zenith angle" ;
		VZA:valid_min = 0.f ;
		VZA:valid_max = 55.f ;
	float air_pressure(air_pressure) ;
		air_pressure:long_name = "Surface pressure" ;
		air_pressure:units = "hPa" ;
		air_pressure:valid_min = 800.f ;
		air_pressure:valid_max = 1030.f ;
		air_pressure:standard_name = "air_pressure_at_sea_level" ;
	float water_vapour(water_vapour) ;
		water_vapour:long_name = "Total column water vapour" ;
		water_vapour:units = "g cm-2" ;
		water_vapour:valid_min = 0.f ;
		water_vapour:valid_max = 5.f ;
	int AMIN(AMIN) ;
		AMIN:long_name = "Aerosol model index number" ;
		AMIN:valid_min = 1 ;
		AMIN:valid_max = 40 ;
	float T550(T550) ;
		T550:long_name = "Aerosol optical thickness" ;
		T550:valid_min = 0.f ;
		T550:valid_max = 4.f ;
		T550:standard_name = "atmosphere_optical_thickness_due_to_aerosol" ;
	int channel(channel) ;
		channel:long_name = "Channel index number" ;
		channel:valid_min = 1 ;
		channel:valid_max = 4 ;
	uc VGT_R_atm(ADA, SZA, VZA, air_pressure, water_vap., T550, AMIN, channel) ;
		VGT_R_atm:long_name = "Atmospheric scattering term" ;
		VGT_R_atm:scale_factor = 0.004;
		VGT_R_atm:valid_min = 0 ;
		VGT_R_atm:valid_max = 250 ;
	float t(SZA, air_pressure, water_vapour, T550, AMIN, channel) ;
		t:long_name = "Atmospheric transmission" ;
		t:valid_min = 0.0 ;
		t:valid_max = 1.0 ;
	float rho_atm(air_pressure, water_vapour, T550,  AMIN, channel) ;
		rho_atm:long_name = "Atmospheric bihemispherical Albedo" ;
		rho_atm:valid_min = 0.0 ;
		rho_atm:valid_max = 1.0 ;
	float C_O3(channel) ;
		C_O3:long_name = "Ozone correction factor" ;
		C_O3:valid_min = 0.0 ;
		C_O3:valid_max = 1.0 ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "VGT S radiative transfer simulation dataset" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-L2-SD-08-S-BC-IODD" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "S3__SY_2_VSRTAX_20101201T000000_20110301T000000_20101207T120000__BC__D_NT_AUX_01.nc" ;
		:creation_time = "20101207T120000Z" ;
		:validity_start = "20101201T000000Z" ;
		:validity_stop = "20110301T000000Z" ;
data:

 ADA = 0, 6, 12, 18, 24, 30, 36, 42, 48, 54, 60, 66, 72, 78, 84, 90, 96, 102, 
    108, 114, 120, 126, 132, 138, 144, 150, 156, 162, 168, 174, 180 ;

 air_pressure = 800, 900, 1000, 1030 ;

 water_vapour = 0.0, 2.0, 5.0 ;

 T550 = 0, 0.05, 0.1, 0.2, 0.4, 0.6, 1, 1.5, 2, 3, 4 ;
 
 channel = 1, 2, 3, 4 ;

}