netcdf S3__SY_2_VPSRAX_20120101T000000_20140101T000000_20120101T000000__BC__D_NT_AUX_00 {
dimensions:
    wavelength = 914 ;

variables:
    float wavelength(wavelength) ;
        wavelength:units = "nm" ;
        wavelength:valid_min = 410.0 ;
        wavelength:valid_max = 1800.0 ;
    float B0_SRF(wavelength) ;
        B0_SRF:valid_min = 0.0 ;
        B0_SRF:valid_max = 1.0 ;
    float B2_SRF(wavelength) ;
        B2_SRF:valid_min = 0.0 ;
        B2_SRF:valid_max = 1.0 ;
    float B3_SRF(wavelength) ;
        B3_SRF:valid_min = 0.0 ;
        B3_SRF:valid_max = 1.0 ;
    float MIR_SRF(wavelength) ;
        MIR_SRF:valid_min = 0.0 ;
        MIR_SRF:valid_max = 1.0 ;
    float solar_irradiance(wavelength) ;
        solar_irradiance:units = "mW m-2 nm-1";
        solar_irradiance:valid_min = 0.0 ;
        solar_irradiance:valid_max = 10000.0 ;

// global attributes:
        :Conventions = "CF-1.4" ;
        :title = "VGT P spectral response function dataset" ;
        :institution = "Brockmann Consult GmbH" ;
        :source = "TBD" ;
        :history = "" ;
        :comment = "" ;
        :references = "S3-L2-SD-08-S-BC-IODD" ;
        :contact = "info@brockmann-consult.de" ;
        :netCDF_version = "netCDF-4" ;
        :dataset_name = "S3__SY_2_VPSRAX_20120101T000000_20140101T000000_20120101T000000__BC__D_NT_AUX_00.nc" ;
        :creation_time = "20120101T000000Z" ;
        :validity_start = "20140101T000000Z" ;
        :validity_stop = "20120101T000000Z" ;
data:

    wavelength = ${WAVELENGTH} ;

    B0_SRF = ${B0_SRF} ;

    B2_SRF = ${B2_SRF} ;

    B3_SRF = ${B3_SRF} ;

    MIR_SRF = ${MIR_SRF} ;

    solar_irradiance = ${SOLAR_IRRADIANCE} ;
}
