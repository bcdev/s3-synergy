netcdf S3__SY_2_VSRTAX_20120101T000000_20140101T000000_20120101T000000__BC__D_NT_AUX_00 {
dimensions:
    AMIN = 40 ;
    ADA = 31 ;
    SZA = 21 ;
    VZA = 18 ;
    air_pressure = 4 ;
    water_vapour = 3 ;
    T550 = 11 ;
    VGT_channel = 4;
variables:
    float ADA(ADA) ;
        ADA:long_name = "Azimuth difference angle" ;
        ADA:units = "degrees" ;
        ADA:valid_min = 0.f ;
        ADA:valid_max = 180.f ;
    float SZA(SZA) ;
        SZA:long_name = "Solar zenith angle" ;
        SZA:units = "degrees" ;
        SZA:valid_min = 0.f ;
        SZA:valid_max = 70.f ;
        SZA:standard_name = "solar_zenith_angle" ;
    float VZA(VZA) ;
        VZA:long_name = "View zenith angle" ;
        VZA:valid_min = 0.f ;
        VZA:valid_max = 55.f ;
    float air_pressure(air_pressure) ;
        air_pressure:long_name = "Surface pressure" ;
        air_pressure:units = "hPa" ;
        air_pressure:valid_min = 800.f ;
        air_pressure:valid_max = 1030.f ;
        air_pressure:standard_name = "air_pressure_at_sea_level" ;
    float water_vapour(water_vapour) ;
        water_vapour:long_name = "Total column water vapour" ;
        water_vapour:units = "g cm-2" ;
        water_vapour:valid_min = 0.f ;
        water_vapour:valid_max = 5.f ;
    short AMIN(AMIN) ;
        AMIN:long_name = "Aerosol model index number" ;
        AMIN:valid_min = 1 ;
        AMIN:valid_max = 40 ;
    float T550(T550) ;
        T550:long_name = "Aerosol optical thickness" ;
        T550:valid_min = 0.f ;
        T550:valid_max = 4.f ;
        T550:standard_name = "atmosphere_optical_thickness_due_to_aerosol" ;
    short VGT_channel(VGT_channel) ;
        VGT_channel:long_name = "VGT channel index number" ;
        VGT_channel:valid_min = 1 ;
        VGT_channel:valid_max = 4 ;
    ubyte VGT_R_atm(ADA, SZA, VZA, air_pressure, water_vapour, T550, AMIN, VGT_channel) ;
        VGT_R_atm:long_name = "Atmospheric scattering term" ;
        VGT_R_atm:scale_factor = 0.004;
        VGT_R_atm:valid_min = 0 ;
        VGT_R_atm:valid_max = 250 ;
        VGT_R_atm:_DeflateLevel = 9;
    float t(SZA, air_pressure, water_vapour, T550, AMIN, VGT_channel) ;
        t:long_name = "Atmospheric transmission" ;
        t:valid_min = 0.0 ;
        t:valid_max = 1.0 ;
        t:_DeflateLevel = 9;
    float rho_atm(air_pressure, water_vapour, T550,  AMIN, VGT_channel) ;
        rho_atm:long_name = "Atmospheric bihemispherical Albedo" ;
        rho_atm:valid_min = 0.0 ;
        rho_atm:valid_max = 1.0 ;
        rho_atm:_DeflateLevel = 9;
    float C_O3(VGT_channel) ;
        C_O3:long_name = "Ozone correction factor" ;
        C_O3:valid_min = 0.0 ;
        C_O3:valid_max = 1.0 ;

// global attributes:
        :Conventions = "CF-1.4" ;
        :title = "VGT S radiative transfer simulation dataset" ;
        :institution = "Brockmann Consult GmbH" ;
        :source = "" ;
        :history = "" ;
        :comment = "" ;
        :references = "S3-L2-SD-08-S-BC-IODD" ;
        :contact = "info@brockmann-consult.de" ;
        :netCDF_version = "netCDF-4" ;
        :dataset_name = "S3__SY_2_VSRTAX_20120101T000000_20140101T000000_20120101T000000__BC__D_NT_AUX_00.nc" ;
        :creation_time = "20120101T000000Z" ;
        :validity_start = "20140101T000000Z" ;
        :validity_stop = "20120101T000000Z" ;
data:

    ADA = 0.f, 6.f, 12.f, 18.f, 24.f, 30.f, 36.f, 42.f, 48.f, 54.f, 60.f, 66.f, 72.f, 78.f, 84.f, 90.f, 96.f, 102.f,
        108.f, 114.f, 120.f, 126.f, 132.f, 138.f, 144.f, 150.f, 156.f, 162.f, 168.f, 174.f, 180.f ;

    SZA = 0.f, 3.5f, 7.f, 11.5f, 14.f, 17.5f, 21.f, 24.5f, 28.f, 31.5f, 35.f, 38.5f, 42.f, 45.5f, 49.f, 52.5f, 56.f,
        59.5f, 63.f, 66.5f, 70.f ;

    VZA = 0.f, 3.5f, 7.f, 10.5f, 14.f, 17.5f, 21.f, 24.5f, 28.f, 31.f, 34.f, 37.f, 40.f, 43.f, 46.f, 49.f, 52.f, 55.f ;

    air_pressure = 800.f, 900.f, 1000.f, 1030.f ;

    water_vapour = 0.f, 2.f, 5.f ;

    AMIN = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 20, 21, 22, 23,
        24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 38, 39, 40 ;

    T550 = 0.f, 0.05f, 0.1f, 0.2f, 0.4f, 0.6f, 1.f, 1.5f, 2.f, 3.f, 4.f ;

    VGT_channel = 1, 2, 3, 4 ;

    VGT_R_atm = ${VGT_R_ATM} ;

    t  = ${T} ;

    rho_atm  = ${RHO_ATM} ;

    C_O3 =  0.f, 0.f, 0.f, 0.f ;
}