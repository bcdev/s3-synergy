netcdf SLST_NAD_RADIANCE_S${i} {
dimensions:
	N_SCAN_SLST_NAD_05km_L1C = 35200 ;
	N_PIX_SLST_NAD_05km_L1C = 2200 ;
variables:
	short TOA_Radiance_Meas(N_SCAN_SLST_NAD_05km_L1C, N_PIX_SLST_NAD_05km_L1C) ;
		TOA_Radiance_Meas:long_name = "" ;
		TOA_Radiance_Meas:standard_name = "" ;
		TOA_Radiance_Meas:units = "W.m-2.sr-1.um-1" ;
		TOA_Radiance_Meas:add_offset = 0.f ;
		TOA_Radiance_Meas:scale_factor = 1.f ;
		TOA_Radiance_Meas:valid_min = -32767 ;
		TOA_Radiance_Meas:valid_max = 32767 ;
		TOA_Radiance_Meas:_FillValue = -32768s ;
	ubyte exception(N_SCAN_SLST_NAD_05km_L1C, N_PIX_SLST_NAD_05km_L1C) ;
		exception:long_name = "" ;
		exception:standard_name = "" ;
		exception:flag_masks = 1UB, 2UB, 4UB, 8UB, 16UB, 32UB, 64UB, 128UB ;
		exception:flag_meanings = "ISP_absent pixel_absent not_decompressed no_signal saturation invalid_radiance no_parameters unfilled_pixel" ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "SYN L1c test data" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "Sentinel-3 SYN" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-RS-TAF-SY-01247" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:Data_set_name = "SLST_NAD_RADIANCE_S${i}.nc" ;
}
