netcdf s3__sy_2_vpcpax {
dimensions:
	tcl_length = 4 ;
	tsn_length = 5 ;
	tsh_length = 1 ;
variables:
	float tcl(tcl_length) ;
		tcl:long_name = "Thresholds applied for cloud detection" ;
	float tsn(tsn_length) ;
		tcl:long_name = "Thresholds applied for snow/ice detection" ;
	float tsh(tsh_length) ;
		tcl:long_name = "Thresholds applied for cloud shadow detection" ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "SYN L2 configuration parameters dataset" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-L2-SD-08-S-BC-IODD" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "S3__SY_2_VPCPAX_20110701T000000_20120701T000000_20112007T120000__BC__D_NT_AUX_01.nc" ;
		:creation_time = "20110720T120000Z" ;
		:validity_start = "20110701T000000Z" ;
		:validity_stop = "20120701T000000Z" ;

data:

    tcl = 0.2465f, 0.09f, 0.36f, 0.16f ;

    tsn = 0.3075f, 0.2405f, -0.3865f, 0.0435f, 0.0385f ;

    tsh = 0.2f ;
}
