netcdf GEOLOCATION_REF {
dimensions:
	N_LINE_OLC = 60000 ;
	N_DET_CAM = 740 ;
	N_CAM = 5 ;
variables:
	int Geodetic_Latitude(N_CAM, N_LINE_OLC, N_DET_CAM) ;
		Geodetic_Latitude:long_name = "DEM_corrected_geodetic_latitude" ;
		Geodetic_Latitude:units = "degrees_north" ;
		Geodetic_Latitude:valid_min = -90000000 ;
		Geodetic_Latitude:valid_max = 90000000 ;
	int Longitude(N_CAM, N_LINE_OLC, N_DET_CAM) ;
		Longitude:long_name = "DEM_corrected_longitude" ;
		Longitude:units = "degrees_east" ;
		Longitude:valid_min = -180000000 ;
		Longitude:valid_max = 180000000 ;
	short Altitude(N_CAM, N_LINE_OLC, N_DET_CAM) ;
		Altitude:long_name = "DEM_corrected_altitude" ;
		Altitude:units = "m" ;
		Altitude:valid_min = -1000 ;
		Altitude:valid_max = 9000 ;

${Global_Attributes}
}
