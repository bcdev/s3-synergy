netcdf ${CDL_File_Basename} {
dimensions:
	N_DET_SLST_05km = 4 ;
	N_SCAN_SLST_ALT_L1C = 8800 ;
variables:
	double band_centre(N_DET_SLST_05km) ;
		band_centre:long_name = "TBD" ;
		band_centre:standard_name = "radiation_wavelength" ;
		band_centre:units = "m" ;
	double bandwidth(N_DET_SLST_05km) ;
		bandwidth:long_name = "TBD" ;
		bandwidth:standard_name = "TBD" ;
		bandwidth:units = "m" ;
	double solar_irradiance(N_DET_SLST_05km) ;
		solar_irradiance:long_name = "TBD" ;
		solar_irradiance:standard_name = "TBD" ;
		solar_irradiance:units = "W.m-1.um-1" ;

${Global_Attributes}
}
