netcdf vgt_p_auxdata {
dimensions:
	AMIN = 40 ;
	ADA = 10 ;
	SZA = 7 ;
	VZA = 6 ;
	air_pressure = 4 ;
	water_vapour = 3 ;
	T550 = 6 ;
	wavelength = 914;
variables:
	float ADA(ADA) ;
		ADA:long_name = "Azimuth difference angle" ;
		ADA:units = "degrees" ;
		ADA:valid_min = 0.f ;
		ADA:valid_max = 180.f ;
	float SZA(SZA) ;
		SZA:long_name = "Solar zenith angle" ;
		SZA:units = "degrees" ;
		SZA:valid_min = 0.f ;
		SZA:valid_max = 70.f ;
		SZA:standard_name = "solar_zenith_angle" ;
	float VZA(VZA) ;
		VZA:long_name = "View zenith angle" ;
		VZA:valid_min = 0.f ;
		VZA:valid_max = 55.f ;
	float air_pressure(air_pressure) ;
		air_pressure:long_name = "Surface pressure" ;
		air_pressure:units = "hPa" ;
		air_pressure:valid_min = 800.f ;
		air_pressure:valid_max = 1030.f ;
		air_pressure:standard_name = "air_pressure_at_sea_level" ;
	float water_vapour(water_vapour) ;
		water_vapour:long_name = "Total column water vapour" ;
		water_vapour:units = "g cm-2" ;
		water_vapour:valid_min = 0.f ;
		water_vapour:valid_max = 5.f ;
	int AMIN(AMIN) ;
		AMIN:long_name = "Aerosol model index number" ;
		AMIN:valid_min = 1 ;
		AMIN:valid_max = 40 ;
	float T550(T550) ;
		T550:long_name = "Aerosol optical thickness" ;
		T550:valid_min = 0.f ;
		T550:valid_max = 4.f ;
		T550:standard_name = "atmosphere_optical_thickness_due_to_aerosol" ;
	float wavelength(wavelength) ;
		wavelength:long_name = "Wavelength" ;
		wavelength:units = "nm" ;
		wavelength:valid_min = 410.0 ;
		wavelength:valid_max = 1800.0 ;
	uc R_atm(wavelength, T550, water_vapour, air_pressure, VZA, SZA, ADA, AMIN) ;
		R_atm:long_name = "Atmospheric scattering term" ;
		R_atm:scale_factor = 0.004;
		R_atm:valid_min = 0 ;
		R_atm:valid_max = 250 ;
	float t(wavelength, T550, water_vapour, air_pressure, SZA, AMIN) ;
		t:long_name = "Atmospheric transmission" ;
		t:valid_min = 0.0 ;
		t:valid_max = 1.0 ;
	float rho_atm(wavelength, T550, water_vapour, air_pressure, AMIN) ;
		rho_atm:long_name = "Atmospheric bihemispherical Albedo" ;
		rho_atm:valid_min = 0.0 ;
		rho_atm:valid_max = 1.0 ;
	float C_O3(wavelength) ;
		C_O3:long_name = "Ozone correction factor" ;
		C_O3:valid_min = 0.0 ;
		C_O3:valid_max = 1.0 ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "VGT-P auxiliary data" ;
		:institution = "Brockmann Consult" ;	// TBD
		:source = "The method of production of data" ;	// TBD
		:history = "audit trail for modifications of the data" ;	// TBD
		:comment = "??" ;
		:references = "When delivered: reference to ATBD and DPM" ;
		:contact = "{ralf.quast, thomas.storm}@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "vgt_p_auxdata.nc" ;
		:creation_time = "20101130T161206Z" ;
		:validity_start = "???" ;
		:validity_stop = "???" ;
data:

 ADA = 0.0, 18.0, 36.0, 54.0, 72.0, 90.0, 108.0, 126.0, 144.0, 174.0 ;

 air_pressure = 800, 900, 1000, 1030 ;

 water_vapour = 0.0, 2.0, 5.0 ;

 T550 = 0.0, 0.1, 0.4, 1.0, 2.0, 4.0 ;

}