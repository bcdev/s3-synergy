netcdf S3__SY_2_SYCPAX_20120101T000000_20140101T000000_20120101T000000__BC__D_NT_AUX_00 {
dimensions:
	AMIN = 3 ;
	SYN_channel = 30 ;
	OLC_band = 18 ;
	SLS_band = 6 ;
	SLS_view = 2 ;
	NDVI = 4 ;
	NDV_channel = 2 ;
variables:
	short AMIN(AMIN) ;
		AMIN:long_name = "Aerosol model index number" ;
		AMIN:valid_min = 1 ;
		AMIN:valid_max = 40 ;
	short NDV_channel(NDV_channel) ;
		NDV_channel:valid_min = 1 ;
		NDV_channel:valid_max = 30 ;
	short SYN_channel(SYN_channel) ;
		SYN_channel:long_name = "SYN channel index number" ;
		SYN_channel:valid_min = 1 ;
		SYN_channel:valid_max = 30 ;
	short OLC_band(OLC_band) ;
		OLC_band:valid_min = 1 ;
		OLC_band:valid_max = 21 ;
	short SLS_band(SLS_band) ;
		SLS_band:valid_min = 1 ;
		SLS_band:valid_max = 6 ;
	short SLS_view(SLS_view) ;
		SLS_view:valid_min = 1 ;
		SLS_view:valid_max = 2 ;
	float NDVI(NDVI) ;
		NDVI:long_name = "Normalized difference vegetation index" ;
		NDVI:valid_min = -1.0f ;
		NDVI:valid_max = 1.0f ;
	float R_soil(SYN_channel) ;
		R_soil:valid_min = 0.0f ;
		R_soil:valid_max = 1.0f ;
	float R_veg(SYN_channel) ;
		R_veg:valid_min = 0.0f ;
		R_veg:valid_max = 1.0f ;
	float weight_spec(SYN_channel) ;
		weight_spec:valid_min = 0.0f ;
		weight_spec:valid_max = 1.0f ;
	float weight_ang(SLS_view, SLS_band) ;
		weight_ang:valid_min = 0.0f ;
		weight_ang:valid_max = 1.0f ;
	float weight_ang_tot(NDVI) ;
		weight_ang_tot:valid_min = 0.0f ;
		weight_ang_tot:valid_max = 1.0f ;
	float T550_ini ;
		T550_ini:valid_min = 0.0f ;
		T550_ini:valid_max = 0.5f ;
	float v_ini(SLS_view) ;
		v_ini:valid_min = 0.0f ;
		v_ini:valid_max = 1.0f ;
	float w_ini(SLS_band) ;
		v_ini:valid_min = 0.0f ;
		v_ini:valid_max = 1.0f ;
	
	float gamma ;
	float kappa ;
	ubyte ave_square ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "SYN L2 configuration parameters dataset" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-L2-SD-08-S-BC-IODD" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "S3__SY_2_SYCPAX_20120101T000000_20140101T000000_20120101T000000__BC__D_NT_AUX_00.nc" ;
		:creation_time = "20120101T000000Z" ;
		:validity_start = "20140101T000000Z" ;
		:validity_stop = "20120101T000000Z" ;

data:

    AMIN = 1, 2, 3 ;

    NDV_channel = 9, 17 ;

    SYN_channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
        19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30 ;
 
    OLC_band = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 16, 17, 18, 19, 21 ;

    SLS_band = 1, 2, 3, 4, 5, 6 ;

    SLS_view = 1, 2 ;
 
    NDVI = -1.f, 0.1f, 0.7f, 1.f ;

    weight_spec = 1.f, 1.f, 1.f, 1.f, 1.f, 1.f, 1.f, 1.f, 1.f, 1.f, 0.05f, 0.05f, 0.05f, 0.05f, 0.05f, 0.05f, 0.05f, 0.05f, 1.f, 1.f, 0.05f, 0.05f, 1.f, 1.f, 1.f, 1.f, 0.05f, 0.05f, 1.f, 1.f ;
 
    weight_ang = 1.5f, 1.f, 0.5f, 0.5f, 1.f, 1.f, 1.5f, 1.f, 0.5f, 0.5f, 1.f, 1.f;
 
    weight_ang_tot = 1.f, 1.f, 0.5f, 0.5f ;
 
    T550_ini = 0.1f ;
 
    v_ini = 0.5f, 0.3f ;
 
    w_ini = 0.1f, 0.1f, 0.1f, 0.1f, 0.1f, 0.1f ;

    R_soil = ${R_SOIL} ;

    R_veg = ${R_VEG} ;

    gamma = 0.3f ;
 
    kappa = 1.58f ;
  
    ave_square = 8 ;
}
