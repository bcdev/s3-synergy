netcdf ${CDL_File_Basename} {
dimensions:
	N_OLC_L1B_TP = 72226 ;
variables:
	int OLC_L1b_TP_Latitude(N_OLC_L1B_TP) ;
		OLC_L1b_TP_Latitude:long_name = "geodetic_latitude_at_tie_points" ;
		OLC_L1b_TP_Latitude:units = "degrees_north" ;
		OLC_L1b_TP_Latitude:valid_min = -90000000 ;
		OLC_L1b_TP_Latitude:valid_max = 90000000 ;
	int OLC_L1b_TP_Longitude(N_OLC_L1B_TP) ;
		OLC_L1b_TP_Longitude:long_name = "geodetic_longitude_at_tie_points" ;
		OLC_L1b_TP_Longitude:units = "degrees_east" ;
		OLC_L1b_TP_Longitude:valid_min = -180000000 ;
		OLC_L1b_TP_Longitude:valid_max = 180000000 ;
	float sea_level_pressure(N_OLC_L1B_TP) ;
		sea_level_pressure:long_name = "mean_sea_level_pressure" ;
		sea_level_pressure:standard_name = "air_pressure_at_sea_level" ;
		sea_level_pressure:units = "hPa" ;
		sea_level_pressure:valid_min = 0.f ;
		sea_level_pressure:_FillValue = -1.f ;
		sea_level_pressure:coordinates = "OLC_L1b_TP_Latitude OLC_L1b_TP_Longitude" ;
	float total_ozone(N_OLC_L1B_TP) ;
		total_ozone:long_name = "total_columnar_ozone" ;
		total_ozone:standard_name = "atmosphere_mass_content_of_ozone" ;
		total_ozone:units = "kg.m-2" ;
		total_ozone:valid_min = 0.f ;
		total_ozone:_FillValue = -1.f ;
		total_ozone:coordinates = "OLC_L1b_TP_Latitude OLC_L1b_TP_Longitude" ;
	float total_water_vapour(N_OLC_L1B_TP) ;
		total_water_vapour:long_name = "total_columnar_water_vapour" ;
		total_water_vapour:standard_name = "atmosphere_water_vapour_content" ;
		total_water_vapour:units = "g.cm-2" ;
		total_water_vapour:valid_min = 0.f ;
		total_water_vapour:_FillValue = -1.f ;
		total_water_vapour:coordinates = "OLC_L1b_TP_Latitude OLC_L1b_TP_Longitude" ;

${Global_Attributes}
}
