netcdf syn_config_params {
dimensions:
	N_AMIN = TBD ;
	SYN_channel = 30 ;
	NDVI = 4 ;
	NDV_channel_dim = 2 ; // dimension needed for variable 'NDV_channel'
variables:
	int AMIN(N_AMIN) ;
		AMIN:long_name = "Aerosol model index number" ;
		AMIN:valid_min = 1 ;
		AMIN:valid_max = 40 ;
	int NDV_channel(NDV_channel_dim) ;
		NDV_channel:valid_min = 1 ;
		NDV_channel:valid_max = 30 ;
	int SYN_channel(SYN_channel) ;
		SYN_channel:long_name = "SYN channel index number" ;
		SYN_channel:valid_min = 1 ; // IODD says 25, which would clash with the proposed dataset
		SYN_channel:valid_max = 30 ;
	float NDVI(NDVI) ;
		NDVI:long_name = "Normalized difference vegetation index" ;
		NDVI:valid_min = -1.0 ;
		NDVI:valid_max = 1.0 ;
	float R_soil(SYN_channel) ;
		R_soil:valid_min = 0.0 ;
		R_soil:valid_max = 1.0 ;
	float R_veg(SYN_channel) ;
		R_veg:valid_min = 0.0 ;
		R_veg:valid_max = 1.0 ;
	float w(SYN_channel) ;
		w:valid_min = 0.0 ;
		w:valid_max = 1.0 ;
	float angular_weight(NDVI) ;
		angular_weight:valid_min = 0.0 ;
		angular_weight:valid_max = 1.0 ;
	uc averaging_window ;		

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "syn config parameters" ;
		:institution = "Brockmann Consult" ;	// TBD
		:source = "The method of production of data" ;	// TBD
		:history = "audit trail for modifications of the data" ;	// TBD
		:comment = "??" ;
		:references = "When delivered: reference to ATBD and DPM" ;
		:contact = "{ralf.quast, thomas.storm}@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "syn_config_params.nc" ;
		:creation_time = "20101130T161206Z" ;
		:validity_start = "???" ;
		:validity_stop = "???" ;
data:

 NDV_channel = 9, 17 ;

 SYN_channel = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18,
    19, 20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30 ;
 
 NDVI = -1.0, 0.1, 0.7, 1.0 ;

 angular_weight = 1.0, 1.0, 0.5, 0.5 ;

 averaging_window = 8 ;
 
}