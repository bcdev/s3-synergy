netcdf s3__sy_2_vpsrax {
dimensions:
	wavelength = 914 ;

variables:
	float wavelength(wavelength) ;
		wavelength:units = "nm" ;
		wavelength:valid_min = 410.0 ;
		wavelength:valid_max = 1800.0 ;
	float B0_SRF(wavelength) ;
		B0_SRF:valid_min = 0.0 ;
		B0_SRF:valid_max = 1.0 ;
	float B2_SRF(wavelength) ;
		B2_SRF:valid_min = 0.0 ;
		B2_SRF:valid_max = 1.0 ;
	float B3_SRF(wavelength) ;
		B3_SRF:valid_min = 0.0 ;
		B3_SRF:valid_max = 1.0 ;
	float MIR_SRF(wavelength) ;
		MIR_SRF:valid_min = 0.0 ;
		MIR_SRF:valid_max = 1.0 ;
	float solar_irradiance(wavelength) ;
	    solar_irradiance:units = "mW m-2 nm-1";
		solar_irradiance:valid_min = 0.0 ;
		solar_irradiance:valid_max = 10000.0 ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "VGT P spectral response function dataset" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "TBD" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-L2-SD-08-S-BC-IODD" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "S3__SY_2_VPSRAX_20110701T000000_20120701T000000_20112007T120000__BC__D_NT_AUX_01.nc" ;
		:creation_time = "20101207T120000Z" ;
		:validity_start = "20101201T000000Z" ;
		:validity_stop = "20110301T000000Z" ;
data:

 ADA = 0.f, 18.f, 36.f, 54.f, 72.f, 90.f, 108.f, 126.f, 144.f, 162.f, 180.f ;

 SZA = 0.f, 10.f, 20.f, 30.f, 40.f, 50.f, 60.f, 70.f ;

 VZA = 0.f, 9.5f, 19.f, 28.f, 37.f, 46.f, 55.f ;

 air_pressure = 800.f, 900.f, 1000.f, 1030.f ;

 water_vapour = 0.f, 2.f, 5.f ;

 AMIN = 22 ;

 T550 = 0.f, 0.1f, 0.4f, 1.f, 2.f, 4.f ;

 wavelength = ${WAVELENGTH} ;

 B0_SRF = ${B0_SRF} ;

 B2_SRF = ${B2_SRF} ;

 B3_SRF = ${B3_SRF} ;

 MIR_SRF = ${MIR_SRF} ;

 solar_irradiance = ${SOLAR_IRRADIANCE} ;
}
