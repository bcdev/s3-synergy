netcdf olc_radiance_o1 {
dimensions:
	N_LINE_OLC = 5 ; // 60.000 in actual product
	N_DET_CAM = 4 ;
	N_CAM = 1 ;
variables:
	short TOA_Radiance_Meas(N_CAM, N_LINE_OLC, N_DET_CAM) ;
		TOA_Radiance_Meas:long_name = "TOA_radiances_O1" ;
		TOA_Radiance_Meas:standard_name = "toa_upwelling_spectral_radiance" ;
		TOA_Radiance_Meas:units = "mW.m-2.sr-1.nm-1" ;
		TOA_Radiance_Meas:scale_factor = 1;
		TOA_Radiance_Meas:add_offset = 0 ;
		TOA_Radiance_Meas:valid_min = 1 ;
		TOA_Radiance_Meas:valid_max = 65535 ;
		TOA_Radiance_Meas:_FillValue = 0;
	short error_estimates(N_CAM, N_LINE_OLC, N_DET_CAM) ;
		error_estimates:long_name = "TOA_radiances_O1" ;
		error_estimates:units = "mW.m-2.sr-1.nm-1" ;		
		error_estimates:valid_min = 1 ;
		error_estimates:valid_max = 65535 ;
		error_estimates:_FillValue = 0;
		error_estimates:add_offset = 0 ;
		error_estimates:scaling_factor = 1;		
	
// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "SYN L1c dummmy data" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "Sentinel-3 OLCI" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-RS-TAF-SY-01247" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:Data_set_name = "OLC_RADIANCE_O1.nc" ;
		
data:

 TOA_Radiance_Meas = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19;

 error_estimates = 5, 4, 3, 2, 1 ;
	
}