netcdf S3__SY_2_VSCPAX {
dimensions:
    AMIN = 1 ;
    NDV_channel = 2 ;
variables:
    short AMIN(AMIN) ;
        AMIN:long_name = "Aerosol model index number" ;
        AMIN:valid_min = 1 ;
        AMIN:valid_max = 40 ;
    short NDV_channel(NDV_channel) ;
        NDV_channel:valid_min = 1 ;
        NDV_channel:valid_max = 4 ;

// global attributes:
        :Conventions = "CF-1.4" ;
        :title = "VGT S configuration parameter dataset" ;
        :institution = "Brockmann Consult GmbH" ;
        :source = "" ;
        :history = "" ;
        :comment = "" ;
        :references = "S3-L2-SD-08-S-BC-IODD" ;
        :contact = "info@brockmann-consult.de" ;
        :netCDF_version = "netCDF-4" ;
        :dataset_name = "S3__SY_2_VSCPAX_${VALIDITY_START}_${VALIDITY_STOP}_${CREATION_TIME}__BC__D_NT_AUX_${VERSION}.nc" ;
        :creation_time = "${CREATION_TIME}Z" ;
        :validity_start = "${VALIDITY_START}Z" ;
        :validity_stop = "${VALIDITY_STOP}Z" ;
data:

    AMIN = 1 ;

    NDV_channel = 2, 3 ;
}