netcdf TIME_STAMP_OLC {
dimensions:
	N_LINE_OLC = 60000 ;
variables:
	int64 OLCI_time_stamps(N_LINE_OLC) ;
		OLCI_time_stamps:long_name = "elapsed UTC time since 01 JAN 2000 0h" ;
		OLCI_time_stamps:standard_name = "time" ;
		OLCI_time_stamps:units = "microseconds since 2000-01-01 0:0:0" ;
		OLCI_time_stamps:valid_min = 400000000000000L ;
		OLCI_time_stamps:valid_max = 2000000000000000L ;
		OLCI_time_stamps:_FillValue = -1L ;

${Global_Attributes}
}
