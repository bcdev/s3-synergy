netcdf S3__SY_2_VPRTAX {
dimensions:
    AMIN = 1 ;
    ADA = 11 ;
    SZA = 8 ;
    VZA = 7 ;
    air_pressure = 4 ;
    water_vapour = 3 ;
    T550 = 6 ;
    wavelength = 833;
variables:
    float ADA(ADA) ;
        ADA:long_name = "Azimuth difference angle" ;
        ADA:units = "degrees" ;
        ADA:valid_min = 0.f ;
        ADA:valid_max = 180.f ;
    float SZA(SZA) ;
        SZA:long_name = "Solar zenith angle" ;
        SZA:units = "degrees" ;
        SZA:valid_min = 0.f ;
        SZA:valid_max = 70.f ;
        SZA:standard_name = "solar_zenith_angle" ;
    float VZA(VZA) ;
        VZA:long_name = "View zenith angle" ;
        VZA:valid_min = 0.f ;
        VZA:valid_max = 60.f ;
    float air_pressure(air_pressure) ;
        air_pressure:long_name = "Surface pressure" ;
        air_pressure:units = "hPa" ;
        air_pressure:valid_min = 800.f ;
        air_pressure:valid_max = 1030.f ;
        air_pressure:standard_name = "air_pressure_at_sea_level" ;
    float water_vapour(water_vapour) ;
        water_vapour:long_name = "Total column water vapour" ;
        water_vapour:units = "g cm-2" ;
        water_vapour:valid_min = 0.f ;
        water_vapour:valid_max = 5.f ;
    short AMIN(AMIN) ;
        AMIN:long_name = "Aerosol model index number" ;
        AMIN:valid_min = 1 ;
        AMIN:valid_max = 1 ;
    float T550(T550) ;
        T550:long_name = "Aerosol optical thickness" ;
        T550:valid_min = 0.f ;
        T550:valid_max = 4.f ;
        T550:standard_name = "atmosphere_optical_thickness_due_to_aerosol" ;
    float wavelength(wavelength) ;
        wavelength:long_name = "Wavelength" ;
        wavelength:units = "nm" ;
        wavelength:valid_min = 410.f ;
        wavelength:valid_max = 1800.f ;
    ubyte R_atm(ADA, SZA, VZA, air_pressure, water_vapour, T550, AMIN, wavelength) ;
        R_atm:long_name = "Atmospheric scattering term" ;
        R_atm:scale_factor = 0.004;
        R_atm:valid_min = 0 ;
        R_atm:valid_max = 250 ;
        R_atm:_DeflateLevel = 9;
    float t(SZA, air_pressure, water_vapour, T550, AMIN, wavelength) ;
        t:long_name = "Atmospheric transmission" ;
        t:valid_min = 0.f ;
        t:valid_max = 1.f ;
        t:_DeflateLevel = 9;
    float rho_atm(air_pressure, water_vapour, T550, AMIN, wavelength) ;
        rho_atm:long_name = "Atmospheric bihemispherical Albedo" ;
        rho_atm:valid_min = 0.f ;
        rho_atm:valid_max = 1.f ;
        rho_atm:_DeflateLevel = 9;
    float C_O3(wavelength) ;
        C_O3:long_name = "Ozone correction factor" ;
        C_O3:valid_min = 0.f ;
        C_O3:valid_max = 1.f ;

// global attributes:
        :Conventions = "CF-1.4" ;
        :title = "SYN L2 radiative transfer simulation dataset" ;
        :institution = "Brockmann Consult GmbH" ;
        :source = "" ;
        :history = "" ;
        :comment = "" ;
        :references = "S3-L2-SD-08-S-BC-IODD" ;
        :contact = "info@brockmann-consult.de" ;
        :netCDF_version = "netCDF-4" ;
        :dataset_name = "S3__SY_2_VPRTAX_${VALIDITY_START}_${VALIDITY_STOP}_${CREATION_TIME}__BC__D_NT_AUX_${VERSION}.nc" ;
        :creation_time = "${CREATION_TIME}Z" ;
        :validity_start = "${VALIDITY_START}Z" ;
        :validity_stop = "${VALIDITY_STOP}Z" ;
data:

    ADA = 0.f, 18.f, 36.f, 54.f, 72.f, 90.f, 108.f, 126.f, 144.f, 162.f, 180.f ;

    SZA = 0.f, 10.f, 20.f, 30.f, 40.f, 50.f, 60.f, 70.f ;

    VZA = 0.f, 10.f, 20.f, 30.f, 40.f, 50.f, 60.f ;

    air_pressure = 800.f, 900.f, 1000.f, 1030.f ;

    water_vapour = 0.f, 2.f, 5.f ;
 
    AMIN = 1 ;

    T550 = 0.f, 0.1f, 0.4f, 1.f, 2.f, 4.f ;
 
    wavelength = ${WAVELENGTH} ;

    R_atm = ${R_ATM} ;

    t = ${T} ;

    rho_atm = ${RHO_ATM} ;

    C_O3 = ${C_O3};
}