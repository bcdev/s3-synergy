netcdf S3__SY_2_VPCPAX {
dimensions:
    tcl_length = 4 ;
    tsn_length = 5 ;
    tsh_length = 1 ;
variables:
    float tcl(tcl_length) ;
        tcl:long_name = "Thresholds applied for cloud detection" ;
    float tsn(tsn_length) ;
        tcl:long_name = "Thresholds applied for snow/ice detection" ;
    float tsh(tsh_length) ;
        tcl:long_name = "Thresholds applied for cloud shadow detection" ;

// global attributes:
        :Conventions = "CF-1.4" ;
        :title = "SYN L2 configuration parameters dataset" ;
        :institution = "Brockmann Consult GmbH" ;
        :source = "" ;
        :history = "" ;
        :comment = "" ;
        :references = "S3-L2-SD-08-S-BC-IODD" ;
        :contact = "info@brockmann-consult.de" ;
        :netCDF_version = "netCDF-4" ;
        :dataset_name = "S3__SY_2_VPCPAX_${VALIDITY_START}_${VALIDITY_STOP}_${CREATION_TIME}__BC__D_NT_AUX_${VERSION}.nc" ;
        :creation_time = "${CREATION_TIME}Z" ;
        :validity_start = "${VALIDITY_START}Z" ;
        :validity_stop = "${VALIDITY_STOP}Z" ;

data:

    tcl = 0.2465f, 0.09f, 0.36f, 0.16f ;

    tsn = 0.3075f, 0.2405f, -0.3865f, 0.0435f, 0.0385f ;

    tsh = 0.2f ;
}
