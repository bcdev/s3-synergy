netcdf dataset {
dimensions:
	NDV_channel = 2 ; // dimension needed for variable 'NDV_channel'
variables:
	int NDV_channel(NDV_channel) ;
		NDV_channel:valid_min = 1 ;
		NDV_channel:valid_max = 4 ;

// global attributes:
		:Conventions = "CF-1.4" ;
		:title = "VGT S configuration parameter dataset" ;
		:institution = "Brockmann Consult GmbH" ;
		:source = "" ;
		:history = "" ;
		:comment = "" ;
		:references = "S3-L2-SD-08-S-BC-IODD" ;
		:contact = "info@brockmann-consult.de" ;
		:netCDF_version = "netCDF-4" ;
		:dataset_name = "S3__SY_2_VSCPAX_20101201T000000_20110301T000000_20101207T120000__BC__D_NT_AUX_01.nc" ;
		:creation_time = "20101207T120000Z" ;
		:validity_start = "20101201T000000Z" ;
		:validity_stop = "20110301T000000Z" ;
data:

 NDV_channel = 2, 3 ;
 
}